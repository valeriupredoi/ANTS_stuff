dimensions:
	latitude = 3 ;
	longitude = 4 ;
variables:
	int m01s01i001(latitude, longitude) ;
		m01s01i001:_FillValue = -99 ;
		m01s01i001:um_stash_source = "m01s01i001" ;
		m01s01i001:grid_mapping = "latitude_longitude" ;
	int latitude_longitude ;
		latitude_longitude:grid_mapping_name = "latitude_longitude" ;
		latitude_longitude:longitude_of_prime_meridian = 0. ;
		latitude_longitude:earth_radius = 6371229. ;
	int latitude(latitude) ;
		latitude:axis = "Y" ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	int longitude(longitude) ;
		longitude:axis = "X" ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;

// global attributes:
		:history = "0001-01-01T00:00:00: program arg1 arg2" ;
		:Conventions = "CF-1.7" ;
}
